-- Created by: Peter KURNEV
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BOPDS 

  ---Purpose:  
  -- The package contains classes that implements  
  -- the data structure for  
  -- general fuse and boolean operation algorithms

uses
    MMgt,
    TCollection, 
    TColStd,    
    gp,         
    Bnd,        
    TopAbs,      
    TopoDS, 
    TopTools, 
    IntTools,    
    --    	     
    BOPCol
is 
    --
    -- classes 
    --
    class ShapeInfo; 
    class IndexRange;  
    class DS;  
    class PassKey;   
    class PassKeyBoolean;   
    class PassKeyMapHasher;   
    class Tools;   
    class Iterator;   
    class Pave;    
    class PaveMapHasher;
    class PaveBlock;   
    class CommonBlock;   
    class SubIterator;
    class Point;
    class Curve;
    class FaceInfo; 
    class IteratorSI;
    --
    --  pointers
    --
    pointer PDS to DS from BOPDS;
    pointer PIterator to Iterator from BOPDS;
    pointer PIteratorSI to IteratorSI from BOPDS;
    --
    -- primitives
    --
    imported VectorOfShapeInfo  from BOPDS;
    imported VectorOfIndexRange from BOPDS; 
    imported ListOfPassKeyBoolean from BOPDS; 
    imported ListIteratorOfListOfPassKeyBoolean from BOPDS; 
    imported DataMapOfIntegerListOfInteger from BOPDS; 
    imported MapOfPassKey from BOPDS; 
    imported MapOfPassKeyBoolean from BOPDS; 
    imported VectorOfListOfPassKeyBoolean from BOPDS; 
    imported ListOfPave from BOPDS; 
    imported ListOfPaveBlock from BOPDS; 
    imported VectorOfListOfPaveBlock from BOPDS; 
    imported DataMapOfPaveBlockListOfPaveBlock from BOPDS; 
    imported MapOfPaveBlock from BOPDS; 
    imported DataMapOfPaveBlockListOfInteger from BOPDS; 
    imported DataMapOfPassKeyListOfPaveBlock from BOPDS; 
    imported CoupleOfPaveBlocks from BOPDS; 
    imported DataMapOfShapeCoupleOfPaveBlocks from BOPDS; 
    imported MapOfCommonBlock from BOPDS; 
    imported VectorOfFaceInfo from BOPDS;  
    imported MapOfPave from BOPDS;
    imported IndexedDataMapOfPaveBlockListOfPaveBlock from BOPDS;
    imported DataMapOfIntegerListOfPaveBlock from BOPDS; 
    imported DataMapOfIntegerMapOfPaveBlock from BOPDS;
    imported IndexedMapOfPaveBlock from BOPDS;
    imported IndexedDataMapOfPaveBlockListOfInteger from BOPDS;
    imported IndexedDataMapOfShapeCoupleOfPaveBlocks from BOPDS;
    imported DataMapOfPaveBlockCommonBlock from BOPDS;
    --  
    imported Interf   from BOPDS;   
    imported InterfVV from BOPDS;   
    imported InterfVE from BOPDS;   
    imported InterfVF from BOPDS;   
    imported InterfEE from BOPDS;   
    imported InterfEF from BOPDS;   
    imported InterfFF from BOPDS; 
    imported InterfVZ from BOPDS;  
    imported InterfEZ from BOPDS;  
    imported InterfFZ from BOPDS;  
    imported InterfZZ from BOPDS;  
    --
    imported VectorOfInterfVV from BOPDS; 
    imported VectorOfInterfVE from BOPDS; 
    imported VectorOfInterfVF from BOPDS; 
    imported VectorOfInterfEE from BOPDS; 
    imported VectorOfInterfEF from BOPDS; 
    imported VectorOfInterfFF from BOPDS;  
    imported VectorOfInterfVZ from BOPDS; 
    imported VectorOfInterfEZ from BOPDS; 
    imported VectorOfInterfFZ from BOPDS; 
    imported VectorOfInterfZZ from BOPDS; 
    --  
    imported VectorOfPoint from BOPDS; 
    imported VectorOfCurve from BOPDS; 
    imported VectorOfPave  from BOPDS; 
    --
end BOPDS;

